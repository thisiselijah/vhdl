library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use IEEE.STD_LOGIC_ARITH.ALL;
use IEEE.STD_LOGIC_UNSIGNED.ALL;

entity bird_control is
    Port ( clk : in STD_LOGIC;
           game_state : in std_logic_vector(1 downto 0);
           button : in STD_LOGIC; -- Input for button press
           bird_pos : out INTEGER range 0 to 14);
end bird_control;

architecture Behavioral of bird_control is
    signal bird_y : INTEGER range 0 to 14 := 7; -- Initial position
    signal en, reset : std_logic;
    signal slow_clk : std_logic;
    signal clk_counter : integer := 0;
     
begin
	en <= '1' when game_state = "10";
	
    process(clk, button)
    begin
        if rising_edge(clk) then
			if en = '1' then
				if button = '1' then
					-- Move bird up
					if bird_y > 0 then
						bird_y <= bird_y - 1;
					end if;
				end if;
				-- Gravity effect: bird moves down
				if bird_y < 14 then
					bird_y <= bird_y + 1;
				end if;
			end if;
        end if;
    end process;
    
    bird_pos <= bird_y;
end Behavioral;
