library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
--The state machine
entity game_controller is
    Port ( clk : in STD_LOGIC;
           reset : in STD_LOGIC;
           start_button : in STD_LOGIC;
           collision : in STD_LOGIC;
           bird_x_pos : in INTEGER range 0 to 15; -- Bird's x position
           pipe_pos : in STD_LOGIC_VECTOR(15 downto 0); -- Pipe positions
           game_state : out STD_LOGIC_VECTOR(1 downto 0);
           score : out INTEGER range 0 to 99); -- Player's score
end game_controller;

architecture Behavioral of game_controller is
    type state_type is (WAIT_STATE, START, RUNNING, GAME_OVER);
    signal current_state, next_state : state_type;
    signal internal_score : INTEGER range 0 to 99 := 0; -- Internal score signal
begin
    process(clk, reset)
    begin
        if reset = '1' then
            current_state <= WAIT_STATE;
            internal_score <= 0;
        elsif rising_edge(clk) then
            current_state <= next_state;
            if current_state = RUNNING and bird_x_pos = 2 and pipe_pos(0) = '0' then -- Detect pipe crossing
                if internal_score < 99 then
                    internal_score <= internal_score + 1;
                end if;
            end if;
        end if;
    end process;

    process(current_state, collision, start_button, reset)
    begin
        case current_state is
            when WAIT_STATE =>
                if start_button = '1' then
                    next_state <= START; 
                else
                    next_state <= WAIT_STATE;
                end if;
            when START =>
                if start_button = '1' then
                    next_state <= RUNNING;
                else
                    next_state <= START;
                end if;
            when RUNNING =>
                if collision = '1' then
                    next_state <= GAME_OVER;
                else
                    next_state <= RUNNING;
                end if;
            when GAME_OVER =>
                next_state <= WAIT_STATE; 
        end case;
    end process;

    process(current_state)
    begin
        case current_state is
            when WAIT_STATE   => game_state <= "00";
            when START => game_state <= "01";
            when RUNNING    => game_state <= "10";
            when GAME_OVER  => game_state <= "11";
        end case;
    end process;
    score <= internal_score;
end Behavioral;
